// Substitutes Xilinx IP core for simulation purposes
module clk_wiz_1(output clk_out, input clk_in);
   assign clk_out = clk_in;
endmodule
